module top_module (
    input clk,
    input reset,
    input [7:0] d,
    output [7:0] q
);
  // 0x34 is hexadecimal which is equivalent to 8'h34. as 4 binary bits are required for 1 hexadecimal number.
    always @(negedge clk) begin
        if (reset) q<=8'h34;
        else q <= d;
    end   

endmodule
