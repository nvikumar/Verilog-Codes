module top_module( 
    input [2:0] in,
    output [1:0] out );

  // m = 1: using addition operator
    assign out = in[0] + in[1] + in[2];
    
  // m = 2 : using loop procedural block
    /*
    always @(*) begin
        out = 0;
        for (integer i = 0; i< $bits(in); i = i+1) 
              out = out + in[i];
    end
    */

  // m = 3 : using loop procedural block another method
    /*
    always @(*) begin
        out = 0;
        for (integer i = 0; i< $bits(in); i = i+1) 
              if (in[i])
                  out = out + 1'b1;
    end
    */

  // m = 4 : using truth table - 1
  /*
  // This is a function of 3 inputs. One method is to use a 8-entry truth table:
	// in[2:0] out[1:0]
	// 000      00
	// 001      01
	// 010      01
	// 011      10
	// 100      01
	// 101      10
	// 110      10
	// 111      11
	assign out[0] = (~in[2] & ~in[1] & in[0]) | (~in[2] & in[1] & ~in[0]) | (in[2] & ~in[1] & ~in[0]) | (in[2] & in[1] & in[0]);
	assign out[1] = (in[1] & in[0]) | (in[2] & in[0]) | (in[2] & in[1]);
  */

  // m = 5 : using truth table - 2
  // Yet another method uses behavioural code inside a procedure (combinational always block)
	// to directly implement the truth table:
	/*
	always @(*) begin
		case (in)
			3'd0: out = 2'd0;
			3'd1: out = 2'd1;
			3'd2: out = 2'd1;
			3'd3: out = 2'd2;
			3'd4: out = 2'd1;
			3'd5: out = 2'd2;
			3'd6: out = 2'd2;
			3'd7: out = 2'd3;
		endcase
	end
	*/

endmodule
